library verilog;
use verilog.vl_types.all;
entity testCode_tb is
end testCode_tb;
