library verilog;
use verilog.vl_types.all;
entity yima38_tb is
end yima38_tb;
