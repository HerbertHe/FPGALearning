library verilog;
use verilog.vl_types.all;
entity jishuqi_tb is
end jishuqi_tb;
